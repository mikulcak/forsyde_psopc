-------------------------------------------------------
--! @file
--! @brief The standard top level VHDL file used by the projects after it has been adapted by prepare_vhdl::prepare_vhdl_file()
-------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--! A debouncer is used to connect the board buttons to the VHDL signals
ENTITY debounce IS
  GENERIC(
    counter_size  :  INTEGER := 19); --counter size (19 bits gives 10.5ms with 50MHz clock)
  PORT(
    clk     : IN  STD_LOGIC;  --input clock
    button  : IN  STD_LOGIC;  --input signal to be debounced
    result  : OUT STD_LOGIC); --debounced signal
END debounce;

ARCHITECTURE logic OF debounce IS
  SIGNAL flipflops   : STD_LOGIC_VECTOR(1 DOWNTO 0); --input flip flops
  SIGNAL counter_set : STD_LOGIC;                    --sync reset to zero
  SIGNAL counter_out : STD_LOGIC_VECTOR(counter_size DOWNTO 0) := (OTHERS => '0'); --counter output
BEGIN

  counter_set <= flipflops(0) xor flipflops(1);   --determine when to start/reset counter
  
  PROCESS(clk)
  BEGIN
    IF(clk'EVENT and clk = '1') THEN
      flipflops(0) <= button;
      flipflops(1) <= flipflops(0);
      If(counter_set = '1') THEN                  --reset counter because input is changing
        counter_out <= (OTHERS => '0');
      ELSIF(counter_out(counter_size) = '0') THEN --stable input time is not yet met
        counter_out <= counter_out + 1;
      ELSE                                        --stable input time is met
        result <= flipflops(1);
      END IF;    
    END IF;
  END PROCESS;
END logic;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--! @brief This entity is the top level instantiating all modules.
--! @details The SOPC Builder-generated system and the debouncer (for the reset key) components are instantiated and connected using signals.
--! Additionally, the rightmost green LED is connected to always light up, thereby signalling the success of the FPGA programming.
entity top_level_entity is
	port (
		CLOCK_50 : in std_logic;
		KEY 	: in std_logic_vector(3 downto 0);
		LEDG : out std_logic_vector(8 downto 0);
		LEDR : out std_logic_vector(17 downto 0);
		HEX0 : out std_logic_vector(6 downto 0);
		HEX1 : out std_logic_vector(6 downto 0);
		HEX2 : out std_logic_vector(6 downto 0);
		HEX3 : out std_logic_vector(6 downto 0);
		HEX4 : out std_logic_vector(6 downto 0);
		HEX5 : out std_logic_vector(6 downto 0);
		HEX6 : out std_logic_vector(6 downto 0);
		HEX7 : out std_logic_vector(6 downto 0);
		SRAM_DQ : inout std_logic_vector(15 downto 0);
		SRAM_ADDR : out std_logic_vector(19 downto 0);
		SRAM_UB_N : out std_logic;
		SRAM_LB_N : out std_logic;
		SRAM_CE_N : out std_logic;
		SRAM_OE_N : out std_logic;
		SRAM_WE_N : out std_logic
	);
end top_level_entity;

architecture rtl of top_level_entity is

	component sopc_system is
		port (
			signal clock_0	: in std_logic;
			signal reset_n : in std_logic;
			-- signal out_port_from_the_LEDs_green : out std_logic_vector(7 downto 0)
			-- the_sram
			signal SRAM_ADDR_from_the_sram : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
			signal SRAM_CE_N_from_the_sram : OUT STD_LOGIC;
			signal SRAM_DQ_to_and_from_the_sram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			signal SRAM_LB_N_from_the_sram : OUT STD_LOGIC;
			signal SRAM_OE_N_from_the_sram : OUT STD_LOGIC;
			signal SRAM_UB_N_from_the_sram : OUT STD_LOGIC;
			signal SRAM_WE_N_from_the_sram : OUT STD_LOGIC
		);
	end component sopc_system;

	component debounce is
	generic(
		counter_size  :  INTEGER := 19); --counter size (19 bits gives 10.5ms with 50MHz clock)
	port(
	    clk     : IN  STD_LOGIC;  --input clock
	    button  : IN  STD_LOGIC;  --input signal to be debounced
	    result  : OUT STD_LOGIC 	--debounced signal 
	);
	end component debounce;

	-- signal right_green_led_row : std_logic_vector(7 downto 0) := (others => '0');

	signal debounced_reset_key : std_logic := '0';
	
begin

	-- turn the single LED 8 on to show that the programming worked
	LEDG(8) <= '1';

	-- turn all other LEDs and the seven-segment displays off
	LEDG(7 downto 1) <= (others => '0');

	-- the rightmost green LED shows whether the reset key is pressed
	LEDG(0) <= not debounced_reset_key;
	
	LEDR <= (others => '0');

	HEX7 <= (others => '1');
	HEX6 <= (others => '1');
	HEX5 <= (others => '1');
	HEX4 <= (others => '1');

	HEX3 <= (others => '1');
	HEX2 <= (others => '1');
	HEX1 <= (others => '1');
	HEX0 <= (others => '1');

	reset_key_debounce : debounce
	port map(
		clk => CLOCK_50,
		button => KEY(0),
		result => debounced_reset_key
	);

	-- Instantiate the Nios II system entity generated by the SOPC Builder.
	sopc_system_instance : sopc_system
	port map(
      SRAM_ADDR_from_the_sram => SRAM_ADDR,
      SRAM_CE_N_from_the_sram => SRAM_CE_N,
      SRAM_DQ_to_and_from_the_sram => SRAM_DQ,
      SRAM_LB_N_from_the_sram => SRAM_LB_N,
      SRAM_OE_N_from_the_sram => SRAM_OE_N,
      SRAM_UB_N_from_the_sram => SRAM_UB_N,
      SRAM_WE_N_from_the_sram => SRAM_WE_N,
		-- out_port_from_the_LEDs_green => right_green_led_row,
		clock_0 => CLOCK_50,
		reset_n => debounced_reset_key
		-- reset_n => '1'
	);
	
end rtl;